library IEEE;
use IEEE.std_logic_1164.all;

entity display_uni is
port(
	res_in: in std_logic_vector(5 downto 0);
	disp_out: out std_logic_vector(7 downto 0));
end display_uni;

architecture disp of display_uni is
begin
		with res_in select
			disp_out <= "01000000" when "000000",--0
			        "01111001" when "000001",--1 
					    "00100100" when "000010",--2
					    "00110000" when "000011",--3
					    "00011001" when "000100",--4
					    "00010010" when "000101",--5
					    "00000010" when "000110",--6
					    "01111000" when "000111",--7
					    "00000000" when "001000",--8
					    "00010000" when "001001",--9
					    "01000000" when "001010",--10
					    "01111001" when "001011",--11
					    "00100100" when "001100",--12
					    "00110000" when "001101",--13
					    "00011001" when "001110",--14
					    "00010010" when "001111",--15
					    "00000010" when "010000",--16
					    "01111000" when "010001",--17
					    "00000000" when "010010",--18
					    "00010000" when "010011",--19
					    "01000000" when "010100",--20
					    "01111001" when "010101",--21
					    "00100100" when "010110",--22
					    "00110000" when "010111",--23
					    "00011001" when "011000",--24
					    "00010010" when "011001",--25
					    "00000010" when "011010",--26
					    "01111000" when "011011",--27
					    "00000000" when "011100",--28
					    "00010000" when "011101",--29
					    "01000000" when "011110",--30
					    "01111001" when "011111",--31
              "00100100" when "100000",--32
			        "00110000" when "100001",--33 
					    "00011001" when "100010",--34
					    "00010010" when "100011",--35
					    "00000010" when "100100",--36
					    "01111000" when "100101",--37
					    "00000000" when "100110",--38
					    "00010000" when "100111",--39
					    "01000000" when "101000",--40
					    "01111001" when "101001",--41
					    "00100100" when "101010",--42
					    "00110000" when "101011",--43
					    "00011001" when "101100",--44
					    "00010010" when "101101",--45
					    "00000010" when "101110",--46
					    "01111000" when "101111",--47
					    "00000000" when "110000",--48
					    "00010000" when "110001",--49
					    "01000000" when "110010",--50
					    "01111001" when "110011",--51
					    "00100100" when "110100",--52
					    "00110000" when "110101",--53
					    "00011001" when "110110",--54
					    "00010010" when "110111",--55
					    "00000010" when "111000",--56
					    "01111000" when "111001",--57
					    "00000000" when "111010",--58
					    "00010000" when "111011",--59
					    "01000000" when others;
                        
end disp;
