library IEEE;
use IEEE.std_logic_1164.all;

entity display_dez is
port(
	res_in: in std_logic_vector(4 downto 0);
	disp_out: out std_logic_vector(7 downto 0));
end display_dez;

architecture disp of display_dez is
begin
		with res_in select
			disp_out <= "11000000" when "00000",--0
			        "11000000" when "00001",--1 
					  "11000000" when "00010",--2
					  "11000000" when "00011",--3
					  "11000000" when "00100",--4
					  "11000000" when "00101",--5
					  "11000000" when "00110",--6
					  "11000000" when "00111",--7
					  "11000000" when "01000",--8
					  "11000000" when "01001",--9
					  "11111001" when "01010",--10
					  "11111001" when "01011",--11
					  "11111001" when "01100",--12
					  "11111001" when "01101",--13
					  "11111001" when "01110",--14
					  "11111001" when "01111",--15
					  "11111001" when "10000",--16
					  "11111001" when "10001",--17
					  "11111001" when "10010",--18
					  "11111001" when "10011",--19
					  "10100100" when "10100",--20
					  "10100100" when "10101",--21
					  "10100100" when "10110",--22
					  "10100100" when "10111",--23
					  "10100100" when "11000",--24
					  "10100100" when "11001",--25
					  "10100100" when "11010",--26
					  "10100100" when "11011",--27
					  "10100100" when "11100",--28
					  "10100100" when "11101",--29
					  "10110000" when "11110",--30
					  "10110000" when "11111";--31

end disp;