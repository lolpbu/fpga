library IEEE;
use IEEE.std_logic_1164.all;

entity display_dez is
port(
	res_in: in std_logic_vector(5 downto 0);
	disp_out: out std_logic_vector(7 downto 0));
end display_uni;

architecture disp of display_dez is
begin
		with res_in select
			disp_out <= "11000000" when "000000",--0
			        "11000000" when "000001",--1 
					    "11000000" when "000010",--2
					    "11000000" when "000011",--3
					    "11000000" when "000100",--4
					    "11000000" when "000101",--5
					    "11000000" when "000110",--6
					    "11000000" when "000111",--7
					    "11000000" when "001000",--8
					    "11000000" when "001001",--9

					    "11111001" when "001010",--10
					    "11111001" when "001011",--11
					    "11111001" when "001100",--12
					    "11111001" when "001101",--13
					    "11111001" when "001110",--14
					    "11111001" when "001111",--15
					    "11111001" when "010000",--16
					    "11111001" when "010001",--17
					    "11111001" when "010010",--18
					    "11111001" when "010011",--19

					    "10100100" when "010100",--20
					    "10100100" when "010101",--21
					    "10100100" when "010110",--22
					    "10100100" when "010111",--23
					    "10100100" when "011000",--24
					    "10100100" when "011001",--25
					    "10100100" when "011010",--26
					    "10100100" when "011011",--27
					    "10100100" when "011100",--28
					    "10100100" when "011101",--29

					    "10110000" when "011110",--30
					    "10110000" when "011111",--31
              "10110000" when "100000",--32
			        "10110000" when "100001",--33 
					    "10110000" when "100010",--34
					    "10110000" when "100011",--35
					    "10110000" when "100100",--36
					    "10110000" when "100101",--37
					    "10110000" when "100110",--38
					    "10110000" when "100111",--39

					    "10011001" when "101000",--40
					    "10011001" when "101001",--41
					    "10011001" when "101010",--42
					    "10011001" when "101011",--43
					    "10011001" when "101100",--44
					    "10011001" when "101101",--45
					    "10011001" when "101110",--46
					    "10011001" when "101111",--47
					    "10011001" when "110000",--48
					    "10011001" when "110001",--49

					    "10010010" when "110010",--50
					    "10010010" when "110011",--51
					    "10010010" when "110100",--52
					    "10010010" when "110101",--53
					    "10010010" when "110110",--54
					    "10010010" when "110111",--55
					    "10010010" when "111000",--56
					    "10010010" when "111001",--57
					    "10010010" when "111010",--58
					    "10010010" when "111011",--59
                        
					    "11000000" when others;
                        
end disp;
